//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_env.sv
// Description : TB Environment
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/04/03
//==============================================================================
`ifndef TB_ENV_SV
    `define TB_ENV_SV

`endif // TB_ENV_SV