//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_pkg.sv
// Description : Testbaench Package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/11/19
//==============================================================================
`ifndef TB_PKG_SV
    `define TB_PKG_SV

package tb_pkg;

endpackage : tb_pkg

`endif // TB_PKG_SV