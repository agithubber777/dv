//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : cmn_macros.svh
// Description : Common macros
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/04/04
//==============================================================================
