//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_test_package.sv
// Description : Test Package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/11/19
//==============================================================================
`ifndef TB_TEST_PACKAGE_SV
    `define TB_TEST_PACKAGE_SV

package tb_test_package;

endpackage : tb_test_package

`endif // TB_TEST_PACKAGE_SV