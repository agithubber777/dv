//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_item_pkg.sv
// Description : Sequence Item Package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/11/19
//==============================================================================
`ifndef TB_ITEM_PKG_SV
    `define TB_ITEM_PKG_SV

package tb_item_pkg;

endpackage : tb_item_pkg

`endif // TB_ITEM_PKG_SV