//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : agent_agent_pkg.sv
// Description : Agent package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/09/23
//==============================================================================
`ifndef AGT_AGENT_PKG_SV
    `define AGT_AGENT_PKG_SV

//  Package: agent_agent_pkg
//
package agt_agent_pkg;
    //  Group : Typedefs

    //  Group : Parameters
    
    //  Group : Include
    `include "agt_agent_common.sv"
    
endpackage: agt_agent_pkg


`endif // AGT_AGENT_PKG_SV