//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : cmn_comparator.sv
// Description : Common comparator
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/03/15
//==============================================================================
`ifndef CMN_COMPARATOR_SV
    `define CMN_COMPARATOR_SV

`endif // CMN_COMPARATOR_SV