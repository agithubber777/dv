//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_coverage_collector.sv
// Description : TB Coverage Collector
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/05/17
//==============================================================================
`ifndef TB_COVERAGE_COLLECTOR_SV
    `define TB_COVERAGE_COLLECTOR_SV

`endif // TB_COVERAGE_COLLECTOR_SV