//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_test_pkg.sv
// Description : TB test package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/09/21
//==============================================================================

package tb_test_pkg;

endpackage : tb_test_pkg