//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_seq_pkg.sv
// Description : Sequence Package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/11/19
//==============================================================================
`ifndef TB_SEQ_PKG_SV
    `define TB_SEQ_PKG_SV

package tb_seq_pkg;

endpackage : tb_seq_pkg

`endif // TB_SEQ_PKG_SV