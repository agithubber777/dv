//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_macros.sv
// Description : TB Macros
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/11/19
//==============================================================================