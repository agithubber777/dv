//==============================================================================
// Copyright (C) 2022 agithubber777
//------------------------------------------------------------------------------
// File        : cmn_base_env.sv
// Description : Common class for environment
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2022/10/27
//==============================================================================
`ifndef CMN_BASE_ENV_SV
    `define CMN_BASE_ENV_SV

`endif // CMN_BASE_ENV_SV