//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : top.sv
// Description : TB top file
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/03/15
//==============================================================================
`ifndef TOP_SV
    `define TOP_SV

module top ();
    
endmodule: top

`endif // TOP_SV