//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_vseq_pkg.sv
// Description : Virtual Sequence Package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/11/19
//==============================================================================
`ifndef TB_VSEQ_PKG_SV
    `define TB_VSEQ_PKG_SV

package tb_vseq_pkg;

endpackage : tb_vseq_pkg

`endif // TB_VSEQ_PKG_SV