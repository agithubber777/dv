//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_env_pkg.sv
// Description : TB Environment package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/03/16
//==============================================================================
`ifndef TB_ENV_PKG_SV
    `define TB_ENV_PKG_SV

package tb_env_pkg;
    
    import tb_env_types_pkg::*;

endpackage : tb_env_pkg

`endif // TB_ENV_PKG_SV