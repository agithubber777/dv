//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_scoreboard.sv
// Description : TB Scoreboard
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/04/03
//==============================================================================
`ifndef TB_SCOREBOARD_SV
    `define TB_SCOREBOARD_SV

`endif // TB_SCOREBOARD_SV