//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_env_types_package.sv
// Description : TB Environment types package
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/03/16
//==============================================================================
`ifndef TB_ENV_TYPES_PKG_SV
    `define TB_ENV_TYPES_PKG_SV

package tb_env_types_pkg;
    import uvm_package::*;

    `include "uvm_macros.svh"
    `include "tb_env_macros.svh"

endpackage : tb_env_types_pkg

`endif // TB_ENV_TYPES_PKG_SV