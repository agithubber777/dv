//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : tb_env_macros.svh
// Description : TB environment macros
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/03/16
//==============================================================================
